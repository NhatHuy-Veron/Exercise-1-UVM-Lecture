// FIFO Driver Class
// This class drives transactions to the DUT

// EXERCISE 1 TASK:
// 1. Add class declaration extending from uvm_driver
// 2. Add `uvm_component_utils macro for factory registration
// 3. Add constructor with name and parent parameters
// 4. Add virtual interface handle (will be used in later exercises)

// Example skeleton:
/*
class fifo_driver extends uvm_driver #(fifo_transaction);
  // Factory registration
  
  // Virtual interface handle
  
  // Constructor
  
endclass
*/