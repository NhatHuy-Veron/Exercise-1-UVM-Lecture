// FIFO Monitor Class
// This class observes activity on the FIFO interface

// EXERCISE 1 TASK:
// 1. Add class declaration extending from uvm_monitor
// 2. Add `uvm_component_utils macro for factory registration
// 3. Add constructor with name and parent parameters
// 4. Add virtual interface handle (will be used in later exercises)
// 5. Add analysis port (will be used in later exercises)

// Example skeleton:
/*
class fifo_monitor extends uvm_monitor;
  // Factory registration
  
  // Virtual interface handle
  
  // Analysis port
  
  // Constructor
  
endclass
*/