// FIFO Base Test Class
// This class creates the environment and starts the test

// EXERCISE 1 TASK:
// 1. Add class declaration extending from uvm_test
// 2. Add `uvm_component_utils macro for factory registration
// 3. Add constructor with name and parent parameters
// 4. Add handle for environment
// 5. Add empty build_phase method (to be implemented in Exercise 2)
// 6. Add empty run_phase method (will be used in later exercises)

// Example skeleton:
/*
class fifo_base_test extends uvm_test;
  // Factory registration
  
  // Environment handle
  
  // Constructor
  
  // Build phase method
  
  // Run phase method
  
endclass
*/