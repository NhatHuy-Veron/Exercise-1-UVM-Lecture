// FIFO Scoreboard Class
// This class checks the correctness of the FIFO functionality

// EXERCISE 1 TASK:
// 1. Add class declaration extending from uvm_scoreboard
// 2. Add `uvm_component_utils macro for factory registration
// 3. Add constructor with name and parent parameters
// 4. Add analysis export (will be used in later exercises)
// 5. Add empty build_phase method (to be implemented in Exercise 2)

// Example skeleton:
/*
class fifo_scoreboard extends uvm_scoreboard;
  // Factory registration
  
  // Analysis export
  
  // Constructor
  
  // Build phase method
  
endclass
*/