// FIFO Agent Class
// This class contains driver, monitor and sequencer

// EXERCISE 1 TASK:
// 1. Add class declaration extending from uvm_agent
// 2. Add `uvm_component_utils macro for factory registration
// 3. Add constructor with name and parent parameters
// 4. Add handles for driver, monitor and sequencer
// 5. Add empty build_phase method (to be implemented in Exercise 2)

// Example skeleton:
/*
class fifo_agent extends uvm_agent;
  // Factory registration
  
  // Component handles
  
  // Constructor
  
  // Build phase method
  
endclass
*/