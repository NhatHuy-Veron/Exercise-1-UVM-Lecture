// FIFO Sequence Class
// This class defines the sequence of transactions to be sent to the DUT

// EXERCISE 1 TASK:
// 1. Add class declaration extending from uvm_sequence
// 2. Add `uvm_object_utils macro for factory registration
// 3. Add constructor
// 4. Add empty body task (will be implemented in later exercises)

// Example skeleton:
/*
class fifo_sequence extends uvm_sequence #(fifo_transaction);
  // Factory registration
  
  // Constructor
  
  // Task: body
  
endclass
*/