// FIFO Transaction Class
// This class represents data transferred to/from the FIFO

// EXERCISE 1 TASK:
// 1. Add class declaration extending from uvm_sequence_item
// 2. Add `uvm_object_utils macro for factory registration
// 3. Add constructor
// 4. Add transaction data fields (wr_en, rd_en, wr_data, rd_data, etc.)

// Example skeleton:
/*
class fifo_transaction extends uvm_sequence_item;
  // Factory registration
  
  // Data members
  
  // Constructor
  
endclass
*/