// FIFO Environment Class
// This class contains the agent and scoreboard

// EXERCISE 1 TASK:
// 1. Add class declaration extending from uvm_env
// 2. Add `uvm_component_utils macro for factory registration
// 3. Add constructor with name and parent parameters
// 4. Add handles for agent and scoreboard
// 5. Add empty build_phase method (to be implemented in Exercise 2)

// Example skeleton:
/*
class fifo_environment extends uvm_env;
  // Factory registration
  
  // Component handles
  
  // Constructor
  
  // Build phase method
  
endclass
*/