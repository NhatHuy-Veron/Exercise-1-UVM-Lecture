`timescale 1ns/100ps
`include "uvm_macros.svh"
package pkg;
  import uvm_pkg::*;

  `include "../model/ahb_environment/ahb_transaction.sv"
  `include "../seq/ahb_sequencer.sv"
  `include "../model/ahb_environment/ahb_driver.sv"
  `include "../model/ahb_environment/ahb_monitor.sv"
  `include "../model/ahb_environment/ahb_agent.sv"
  `include "../model/ahb_environment/ahb_scoreboard.sv"
  `include "../model/ahb_environment/ahb_environment.sv"
  `include "../tests/ahb_base_test.sv"
endpackage: pkg