// FIFO Sequencer Class
// This class controls the sequence of transactions sent to the driver

// EXERCISE 1 TASK:
// 1. Add class declaration extending from uvm_sequencer
// 2. Add `uvm_component_utils macro for factory registration
// 3. Add constructor with name and parent parameters

// Example skeleton:
/*
class fifo_sequencer extends uvm_sequencer #(fifo_transaction);
  // Factory registration
  
  // Constructor
  
endclass
*/