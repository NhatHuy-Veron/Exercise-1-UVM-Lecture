module testbench;

  initial begin
    /** Start the UVM test */
    run_test("ahb_base_test");
  end

endmodule